module butterfly (
	input signed  [15:0] Ar, Br, Cr, Dr,
	input signed  [15:0] Ai, Bi, Ci, Di,
	output signed [15:0] out0r, out1r, out2r, out3r,
	output signed [15:0] out0i, out1i, out2i, out3i
);

	// define parameters for twiddle factor here

	parameter signed [15:0] W0r, W0i, W1r, W1i, W2r, W2i, W3r, W3i, W4r, W4i, W5r, W5i, W6r, W6i, W7r, W7i, W8r, W8i, W9r, W9i;
	W0r = 16'b01_00000000000000; // real(W) = 1.000000000000, imag(W) = 0.000000000000
	W0i = 16'b0;
	W1r = 16'b00_11101100100000; // real(W) = 0.923879532511, imag(W) = -0.382683432365  
	W1i = 16'b11_10011110000010; 
	W2r = 16'b00_10110101000001; // real(W) = 0.707106781187, imag(W) = -0.707106781187
	W2i = 16'b11_01001010111111;  
	W3r = 16'b00_01100001111101; // real(W) = 0.382683432365, imag(W) = -0.923879532511
	W3i = 16'b11_00010011011111;  
	W4r = 16'b00_00000000000000; // real(W) = 0.000000000000, imag(W) = -1.000000000000
	W4i = 16'b10_00000000000000;
	W5r = 16'b11_10011110000010; // real(W) = -0.382683432365, imag(W) = -0.923879532511
	W5i = 16'b11_00010011011111;    
	W6r = 16'b11_01001010111111; // real(W) = -0.707106781187, imag(W) = -0.707106781187
	W6i = 16'b11_01001010111111;  
	W7r = 16'b11_00010011011111; // real(W) = -0.923879532511, imag(W) = -0.382683432365
	W7i = 16'b11_10011110000010; 
	W8r = 16'b10_00000000000000; // real(W) = -1.000000000000, imag(W) = -0.000000000000
	W8i = 16'b00_00000000000000;  
	W9r = 16'b11_00010011011111; // real(W) = -0.923879532511, imag(W) = 0.382683432365
	W9i = 16'b00_01100001111101;  
endmodule 