module butterfly (
	input signed [15:0] Ar, Br, Cr, Dr,
	input signed [15:0] Ai, Bi, Ci, Di,
	input signed [7:0] Wr, Wi, // twiddle factor
	output signed[15:0] out1, out2, out3, out4
);


	always @(A, B, C, D) begin

		


	end




endmodule 