module FFT (
	input clk, rst, 
	input [15:0] din_r,
	input [15:0] din_i,  
	output [32:0] dout
		    );





endmodule